interface intf();

endinterface
program testbench(intf i_intf);
  
endprogram